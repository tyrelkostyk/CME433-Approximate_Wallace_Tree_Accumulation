module eight_bit_wallace_tree();

endmodule
