module eight_bit_wallace_tree(
	input [7:0] A, B,
	output [15:0] S
);

wire [12:0] L_12;
wire [10:0] L_23;

eight_bit_wallace_tree_reduc_layer_1 L1 (
	.A(A),
	.B(B),
	.w16385_in_L2(L_12[12]),
	
	.w1_o(S[0]),
	.w2_o(S[1]),
	.w16385_o(S[14]),
	.w32768_o(S[15]),
	
	.w4_o(L_12[0]),
	.w8_o(L_12[1]),
	.w16_o(L_12[2]),
	.w32_o(L_12[3]),
	.w64_o(L_12[4]),
	.w128_o(L_12[5]),
	.w256_o(L_12[6]),
	.w512_o(L_12[7]),
	.w1024_o(L_12[8]),
	.w2048_o(L_12[9]),
	.w4096_o(L_12[10]),
	.w8192_o(L_12[11])
);


eight_bit_wallace_tree_reduc_layer_2 L2 (
	.A(A[5:0]),
	.B(B[7:2]),
	.w8192_in_L3(L_23[10]),
	
	.w4_in(L_12[0]),
	.w8_in(L_12[1]),
	.w16_in(L_12[2]),
	.w32_in(L_12[3]),
	.w64_in(L_12[4]),
	.w128_in(L_12[5]),
	.w256_in(L_12[6]),
	.w512_in(L_12[7]),
	.w1024_in(L_12[8]),
	.w2048_in(L_12[9]),
	.w4096_in(L_12[10]),
	.w8192_in(L_12[11]),
	
	.w4_o(S[2]),
	.w8192_o(S[13]),
	.w16385_o_L1(L_12[12]),

	.w8_o(L_23[0]),
	.w16_o(L_23[1]),
	.w32_o(L_23[2]),
	.w64_o(L_23[3]),
	.w128_o(L_23[4]),
	.w256_o(L_23[5]),
	.w512_o(L_23[6]),
	.w1024_o(L_23[7]),
	.w2048_o(L_23[8]),
	.w4096_o(L_23[9])	
);


endmodule
